module notg(a,y);
  output y;
  input a;
  not(y,a);
endmodule
